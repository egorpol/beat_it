BZh91AY&SY
�0. �_�Pyc����߰����`�Nm*�;i�����Z�KX"�	�M)��������i6� �4@��LRRi���    �L�i�����a�0  ��T��=�14i�@   �MU�7��Fe!��h@4�""j�HL��i��d M4 <�w���	lp?��R�@d���%�]2�UH>�I%���񚪪��� �JI�ԖL�I��2poɻ����P����7��D��ցkIQ)j�DAr��E`�P�P�'X� �(�)T"�t��X8���-V�X��b)���>[5�a.�~�1!ݕ��*�g|o^�sޯ��r�E�V��~ֵ0�9n�����(ƁP��I���8�F5��*������s-d\�sv2n���1me�Z��:�N�;U�5Dqd���>����\�W��R��(rq�2��哑����WK�<��$� HRPH�����йN�צ����-�y�w=�h�=J��loǖ�~($𞒛�	"��NwЉ=���y��F�	�ZL���� :�}M�w�U�+�ç�ѸEXB��;��$�� �\����`n�����<�'��ʇxS�1�X�>�|�il:s٦���۶��8f\����N�,���,��abl�0�;q�jS�T�ݓ;��L:!�em��-��fd뚩KpӳfTr��#��[96�pr �qҀ��s3e�Rt��N,ٻ�$�I�niF#ȗ/a�x8��xa�C["�칧K_2�)�I��my;.ikiN2Ç}�9r��e�ʛ�TT�+l�ʺS)��8SJ)��)�L�r�n�m(�S�8�q)�taӝ�WTkA#��O���i<�o�FdQ�,����I vGR�~�Np��-�A� v���,]�;C(iE��Z���ӥ�Q�2�p��,�t.�$���h�7x^��d��-��1�x ���ӱi%]փ���G"�,��C0���Z�ae-���wZ�%����Z�l ���x��gGm�g�Ӎ��t�Sfs!�X�)�L���y�JeM�4�St��0p��ޅB��IY��Ôi�<q��50��R��MT��|c+�sxR��Ӽ����ѕ-�k�u֮������6l
0,���J���\X�0��3�::-���*�x"o�UҚ��y��PD�hZPIC�q���Y�t�s�`�D9m�e����8ti�����,��M-�5ŭ���m^BxC���{�r�r�vp�xƛ66q;�wt��M�6�̦���Sf0��o7[��SSKP���ԕU��J��y�b�(q� D�j,:�E�i�5�t�q��Z��196en#�\:�o>N���r��D5K�L��N~�p��	�� DDDD@����G�rI�{"�J�����V��xgdK��[���"PΤ��Qe��c23t���Y�\�].-I���J�)%*"eH]�c�Cj�)5$�S�\N�o�*Wf�xC��7�K�ҧu�T�^(�JH%(��C��_�^�쿟���x�c��n%�H'Ƃb>ʎ����"b���������{�f<[��{�>�z9eZT���	�J�9�WF�,px�/��̨�Ң��/����xۇ�KΥ��`�,@H�݆���ل;!a8RQ���	?�}�rMH���p:D܀��CQ��@�}2!��c�J ����$@ M��Zs[�=N.R��F�K[�[�=�õ���U�X�$@������������Au }�GE!�E�^ܰ� uJ�I`�ץ�)%婽�%�c����~��ȉ�\7�V��̨�ug���܇0��<-�F 32���� �.c��H�R>q�Wo{E
�
�fV�ޤK���)����K�*A��ԻA5c&�|z^"��М�5�0\ԻKIcM�V�7 ��DT������o���D�ā��AP��x��XSc��~=uLT���t�K�ڹ��t�š�̏�vm42z(���|�%6O&���1>o�ai�y��;��W-US�l��:�����Lܙ�����Yc�q  I)�o-��-
iWa�P��v��P2��N�u�I���m�zN뼼��	8:g"50h
�}�&q��7S5@�^@kpA�Ll�U��nJ�P��HGo
��U�(:G\���[���
*N��=hב7�F�Z�g�=p��֡eu������~�Ĩ���g��O��r�̵+���2c�v�$�i�A�;{�K�s�x�	�(�a����:p>��G�s�8�T�^�05�Y��B�w����L�P� C �}��)��N��kD.-p��o�g� ��D� �
�B��w$S�	 ��