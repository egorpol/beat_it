BZh91AY&SYxя� 7ߔRyc����߰���� @ `^|� ��(    	q�Y��(*�Hjy#=�4��F�`� f�&� )(�M�2b�h����db0�`!�M0�!�F��JdBh� �     R�=5=F�4 �4�A�$"4�!=7�S12OP��A��fqEY/�����p2 3
�� ��a�eY����-�"����i^h` V%Ga�	z�I2K�*�H��M.p��E�0��*2Uc�Fۼ�I��7OW�t \j��DP��Yr_!���^�tp�a��ƘF� =Ġ9�)}q"/�QM�P�4��}j��j\[5�R�A4fB�o��>�s�ͨ�86\ֵ�]FL����f�-�i�Wo I�b���k'��T����)�Ґ�(c��r0%�SIv�DX�˪7���Bқ���̜V;�B�P ����ff��P�S�/]���3K.�,͒��2d�U1���!+v� 򮶪'Da���Ý�jY�(iEb��^Zص�%��#nT\n���������T2��4j�
�B�>i�]Q>�Ѐ�1�'1���Ħ�VY���UeL��@����lC+]e5���l��K������뿲�ώ��
��"����[�����g�K�m��k��[��C��y��h��^d�H���b�		C/�}�\@��s�n:pz�~��?�gո~�����K4}�����ȹ�\"�9��tv2�RF1M��-+�#f�!{{Bˈ��j�O#mW�&�3����Q�Rll��5����e%��d��Ku�h�~��)H	�3项~�V��6�*�R.p#v���dwK����ʖTy2 Iw��Zj�BDR3\V��V�r�]�m�P�Ȫ�B����@�y ;�_����c����1�ٔ�-�̯2$�<|+;nF"N�D5$����H��h71� Έq��� _�~��9��ׁ��%�	���Ϗ<��H��0�
A�l�pj�C@Sf]�De[F���Jk�|	�������\ `L�ω�"�t��D��aU��anu̸� q4b��V��,�ue��E�m&:��ʭǦ[�Eij{jd�m��[��D�(�4PMYJ� �ݹ��d g�o`I�BE�� �#�w0�`�	�o������.�1&�K�1�ȍ*W�-2cԓ� �_VE�S�v�j��J"�7�1g��0Q}\�h2�D��$� ����\�d�v�6Wt�j
5c>���'�H����L
+��&"�#��v�O���F�1v��N�E@@��,�((8Uf� ���ѧ���>��ƈ"Y�&�j��n��.j��z�5P]�e蚺#L@Q��N1�b�� �2��Cl�<�(�1=;K�8x����Ԣ+� NW�մ����b�3�w��@C^h6L�FXI�`p�v(Q������_Y�Y^G�A��J��7n,=���O4]�����Lu���6l��.n�Z����,i���_��
����>KR$�o竫hS$�1	N��E�K��aL��!r��eC��`==Q��6N��"�\R�DX�M\3����Ơ+W��ܪ>�]�Ńg-h BL4�\"����)M�P�]�$ٟa�0*nO��W���4�
�,ёL���
��GB��R������0��+{�����[u��;cf�%:v����؍���nÐ��蚺�&J�A��FR$Q{\ٗ��<ō���o���1g�l�5�3�o'�b�§�o;�ml��>���?w�}�'�ë$|�|`��o�`�?�/'�,��rI"���}Am�� ��C���8�'*�e��E�+`��ܠ��4�TnZ�a�|Q��q����9�XD�+x�gP:\���!LͣSf!Б�8}�$�Bi?��>Zv�'�Z�;�&����):`Ovz����Q뇳U�0����è!�=EO����"
�\Y7�e��a�[9zL���t ���/[�jq35
�:pgtև~�uiG[�<�,������F�fb�i�	ܱLM�ϓW������U�e�m{�O*����1���fa�3K-?!��/1c-n�u�3� ELhzy}���K���H�g���YUU��ЖLIZ�9��s(�de�t��~����x��ʢ$�$�I$OXD�A[�_� W��+X��Դ�EU[L�+9X*�|�0��!)"@DB�-,��L��b h��wB)��2�je"e��I(d)��T��%E�%�@R��3�Y��[rP��*�$���
��N=\��~�O�Vx��h;�L�����3���Xϝ^e�v����,�f�V��E^&y��� wtHP��r��KeɻI��T_!��&�F����2���B�X��+?�#	�h[P���O�1�hm�v
`Ctm��_թ�ʺ:�D�x x�}�
���N7"�Y;1H���{�Q�
�a2x2��]���Lb�'�R�=����Z�}��LaB�;�.|[��N%�]����$"�j�9D� ܈���a31bF+I��5��ۚ<tlښ|��`O� �Ҕq�^v�@&�D�yA<*m	!̌��Z@j�4@~��� ���<D�A>���v;V� �� �U,8\�(�=����N�Q� �<
!��#�.Tq;6!���9�,�� Nϑ�㣇I��^c��6;��<:�~�ô��w
�4~ɖ
а�=����- 
޶x�0��m�����""���LR�a��Ƞ�p#a��W2�EX������%�<r ��t��-h�KP�aO�2�n�0+;X�[$��$cA��V��Ӝ;���j���L��_@}&�~j[U	ׇ�n��<�X]�@���9���|�k���)O5)��jI�r`EK�d��٬A��{` �ڸW?:�r�{z�zy�h^Wm%.�4���q�۰b	����0u�G����WB^�YWB$��ҝ���g�n{��l�Cg@@�E4��K�~�0!0� ��$%j�-�i�� ��:Ü�nԄ�n��^� �=X������^�͂(�Fu*�̰��՝u�Fp��;��5�-i��܌C%R>�'D�m�t��K�xv��V&�n�H��<3��O~��� ���=s���s����)�ƌ|�