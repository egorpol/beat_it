BZh91AY&SY���� �߀Py����߰����`� ^� a7��UC3�P
d �e�x"$�� � �0�<LT?J�i⟨�� ��P5<��P`2a4``�Oت���L� di�F���M �OС4��� L�   �& �4d40	�10�"
m24'��D�A�F�DѦ�����K �����("�D����D<.�0�H�`PRG��^I@e�QL�TĂwĨ�13G����ׂ�$���"Ȳ������Ȅ�����  �,��� �$��B��"��� � ��ȣ $��`0�H��H��! H����)���I���E�S���f���Q;�6���Ν��H���HZ�u�h�G��m����1�xGAԛJ���5���H0�H�6��[���)u&��ܶ�;'M�E�$�]kt��hrf��X�x�=xki\sk����[�y�u���󷌶G��H����7O]R6�!¼�rs�#�%����v�ZY��nv6w+q��>m��mӚ��ñAۂ��q���<�rJ'Uh����ØB���\�@SiC]�����ݒ%�����]B�����!�FP�&a�T2��)����+b�qOH`�VHvU]03�l��͹E���@$	11�s�^a�dԴ��ǯ	#j��7NR'>n"�F$L>A�6ź�����.ZnN�n�R��s%NURi���p$+�Ӛ����Q�,%�F�*�FO����R��QT�-S&��lfH�5#6�p��z�l'U6=���A�D�b��������C*�f�֍U�jg�ܿB��s>d6�f��iXJ2�Tƚ�7��3����8'�rZ!A($��Sh��,�.�o�#�p��.��C@`k[G)��x��O������F��6��&�� o`d��$�E�*[b�� �+�{x�vdƢ4үS�����0��s�e���a84|�ت揠����˻tq��N!*b\%S,Y �̘��B��-T;_0�Tsu$~h�/g�[���1M�b�.�`��F�S���@�t-�	��C��:P����@C��0�� ��f[}W�'[J��$HL��f9}�����=��/Y� *�
�a�D��xp�3ʠ�[�|�`�L���[�*��g8T�c���ב��&���t���W� �4�c9N��t�A��.��8Xn)���A,Nt\��Hn@�2} Lzz��8���2�V���K�a|'v0��(���^�p�!�QIB��V<�4v%��޳��	AUve���.�J�3�t#�10o��:6-���^(�����I��ю��⑐;: ��5f �h� ��@n>-��>�p`N�@m/
٥�.�{�&��E��>e|ʔ(� "���H�ES�aBNG���JO��& �
����΁Z���uIpヶ�<��I�v$G؎��N�a�l�\�$DBzA�P��U+ va˙Nf��9y1�*,`ބ�@�
��j	 k���<����yy�:��1X&I=�
l]'�my���L>����f�n�{���п7��΋\R@Í�#n�$tp��*I���������HN�$v��Qqہ[S�Z:��
�3���1c��&��mW��2�uy��O`�s�dI�#�}�|h(�.�l�$]�7�v>b�hK��#��LTL6Ԫ%�p��#�c�o
�_`[A�:�zN��m�;�q�TO��d��a`7��ɛ;��Ы(�I �@<!4RBgr�#��t���H�62�/T��eb�in2�c����U>�ZѳFi�E��q*����0��&Z�a1\񚎈7�(v�YH]��`���J���C0�2̌�.��d�B��k��3�儲ESNɊ�ڼS�ǳ(֟Uw�ʠF-���b\F�W���O8`�����g����(�[A0HI0A�c��1)���n�JWM�c%;Oo��n���o�P�IÆ����z�f�t AH������uO$a�+sl.�D����z�����u���]4ܬX���d�`��Bm�0L }uW ��/Q�;E]�b��d��40^�׎h����j���g�Ej�~i���4�$3�w"��"��]�B�;��Ew�"���];Pr���>�쉇��".��1`��\­X�]���J0��.\� OG�⻎�G"8w�$�8���b;@`&�]k�(��m<��a�}��WI�	�q
�������
e���E�i]N�ywuЈ8(Q(!�R���;�7���������GA�D�IRq�%��s���6cG��:�<>7)�<�ᮞ����9]�.H�_����M�I���@:��9��ҹ ����B�L�ic6�ㆷ�qئ�'9�ã�q939(���ԹQ�cd�^(�P4��B�u͙P�:�2�Ɍ�Y��z�1�ƈQ�x��Qe;���U��A��C1���A� �iB@�!�*,v7�\�sC0�+|��+�k"��Q��K�Ctԋ�/"i����}	6Ba��"�5�;�y-�]�v�^�ˍ��%e� �kO*��T7�ƒ�y�.P������0Bj<������UHfAԳ&"]�B�Q#LHk��(]��f��R�Rt(N�H�?^��8��61��m���PR�;� M�`�2e�
>X��}��kq��X�bؖ͊�h���L��Y]A� �R�R)����� �dR��Q!a!@˨��}��l�µ044Hj��Ͳ<�DB�Ą�F����/�m{�l����:�֟�~5�?x󶺸-`�c�6�0�!2��Z|.�	�}�`�����$aiVv���f���2�Z� �����z�2l��+�7E=��$hv'j|��wn�]{�B��m�o��!�҉���

e�^��>�`4�˅��r� w�-Q1�ͅ��^� �w�h "����́��Yx�2S�6�Ϻ�ھ2��Ŵ�EQZ��lD��P%�"�,X.ݬuVQ�Qn�K��Soð�9� ME.Pl��Lzxm��A�����iޒ>'A�A��a��Q��Ǽ��vΫ�,9|��\ �)�d��X9�<�׏�>9�ܝ���
^&J��~��4>�����!��:�V�����ͬ9�N�@��ʒ�9^>��L:�Mn�*�n:AO^�������Ѳ����H1V��D�eǰ�l��0�$!My. ׂ*)BA������,�f�v�(�}�;���,(�oIk���h��=!��A��'7ќW(�=j!��`�ۼ�d�	i$-��꟫n��^w����3�)�q��C�
=j��N_8�I�d��z���LTղ�5`N����@()���*y��Xvi/=:hCa�P�X��mX�9mP+"�'2zW�p�5�/�i0��\����tž `��i��PS"(�;̌*T� �d�j.�䶫�E��X�h��Q��
!@�!A,;/���ȃ��EÞ���۠7Rl��â�����1�,�2����Bv�� �o�2��ܑN$.�p 