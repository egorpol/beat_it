BZh91AY&SY��� A _�Py����߰����`$�w�ղ�=���m��;�k���:�ڤM���ݙͪڭ�Z˶[5C���m��;2��m��VԦ�efZj��_|     j`R�=@H    h 0�?!�*�M      ��� �R�CL� ɂ`&  T� J�SLF� �# CL�ꧤ��� ��  �   "�� F L'��=�S���ˤ� g��Q@h �!x(���! h���
?�.�b
* ��DDG��PT�!�� f-�=����E� �wUV.ߍfS�k�����.�<?y�L�ϣEi��̤/�����K�.�T�Eeͦu�ˇ#����فLN�C֨��!X�VӇ�MNO�E��)�Dl�4(I�B����Q�,�+Mv�O5a�8�_V��F#������Ra�{��Z�d��j�έ'[H;E���Q���S6�C�,f�݆�G��"s-͗[�Z�٣r�-=�]ѡ�T�����;�uģI�{6�Ԣ;��&Di>�ήҠ�Q�ܮv�lr'�s{2�TwW�#w_IM����0�]�3�-a���s`D.���6%~�~�>:-yW��4��f�q�>�����M�3�T�b��ة띶�\����g�u��]�d�4�OX�q2+'[�H����ΐ�g�)�&}xp�wp��e�����&��e��=���u�*�������L0��5�����k��p�t='�R��:��S�l�[�(�o�ل,ۣ���OB{Y��Q�P��m�	u�|�GJt�斛�ɩ�P�/j
,tv���A�J��:��b%f��b�)�;�sH!!v���X���$���v���5�#����E�{�.��D�c�7m�@@�r}�ϯ-t�+`����yX4F����B���M2P��sR�Q�������(�[xh�y��+�N	�[���[T�j��˘�od���]�5�{]l�����hnꖸŚͺ���=�<Wf	���3y�����0f�By̲iϫas��b����d�vP��RƦ���f��� t��} �)x_r�k�B���q��ɧ_C���� �'e��v$�d3Ð�;cW�$tn����8Ct_�m���KH�k����#k76y2{����	��B��D�Of:)�Fn#�e�L�᣽r�R3���4�aFGm�T��������A�
4[���|����0k�[ �:���E{�BW������O�N�����o$m���.|s�zI�:i�����]��c�AX���^��1�{ Ż�{7c�wRoX�-\7b.Ź�C�����K<b��t�����%��%o����ܽ�v�H��U)t/YH?�4mG$��j��Ն�	��돕����uB����M�)ɬ�^��kHߍ��"H�D��p-޹e�\�~f"5�NZk�w.x�f�F�[���<��E��|�;�V_[F"����f�*W6���� �6�b��j�/�ϸ�&���6m�|��{k�N*Y�8�=���$�s�O5���x��>ߨ��K��Rp~��Y����.K\3m]cͯ"����ENS����as��!Λ��G����D�&�Q�L�*K_�)���f�G蹎!����[��|E�#�ݶ)���g�@����l����5��{�X31C�{]����(�R�`��F�?H��b�J��=񉹰u�c�gϽs�v���Ю��#"QN����s(�u�5|�N�Ԧ������H^n�B�B<�|�i�uPR�!�Ò���W�~я�2�`;�Ϸ�*���)�@��ͰZ��:G!����v4���Q�%~���@�0�fm3�e+pE�hs~��xH��H�C�!:�����h8y�$���F�F^"�_QPK�`�C�y`[�ذ���T�۸^��I^��A&}�a��%�c�)��A�J���}�7��~mQ�ü���-*���0��]�pl�ǽ�s�Ցy�/r��
5�N�����k�I�S�v�9}5��[~!�#��Zo�ݭ���Nk��w���~U�/���e�r��[ �l'�lQ,�fS=����D�2���ٙ)�(Pl��瑛Ő�p?AI*a�O]
�O惲�l_�W�J����rg6�B$H�Gꎚ,��N1P�ju~%Vb�g��H2��cfF�uajm���a�L��喞2��c�,<`a��1���vZ7��k�	�j�϶�<�w2V>�-{�	������Z����	�Kx��@��F�>���/
��A���^S�7��NU/\�_я}�9T6�[$����miCyJ�>��p��-غ�(��h��U��:��SX0w�o��3<����w���f�,�T�__��pO���l�aW�C�p��	�u�l��/y�<8!���jLxOV�G�mu���m�}�)��s�z�Rd5ٵFy��X'��=��z�Ahy���]�f]X���������������"nw�*'E=t# �R_F!s�ޒs��v8��P��ɀ�ЛRR	�ׂ!>D�W�"P��y��ֹĚa����2g���v��s�:?��RV
#����{�|k���e��}�&�W��६�ֹT�����r�����o��t3u�8y�����崗�.a`�j� yn��>z�/�y���	Q�r�eQ����b�u�{���?�݊�/�Que7q�a��������{��n�Y]px�%�^}�֞(u"'�'H+GH���N;[Yޣ�ꋳ��w1V�y�b���N�6`�s�Q�Dl5a�"��m���ς 6!5����j����=��)�;=��
�[�(�:ũ`5u�s`��!3D���=��*oA_�Zľ:ٱw��$Y����$�~.��x�QE[��KB�U~b�b`CީfmUQ���k�Ȧ�O�g���d=�����Ņm�a�J���/�q�M��۱�8��,t��E�]��Ī�������S{����k<�kڌ���L���N{4��s�h6�X;Y9�<,����n�(,�C�ǳE�'0��I"������U.������&D��hIX��(o������mK����8�
����S�\�[�A:ua,5��#T�&���o"nn_�'jb��҅_�!F?��&���l-��?z�@��͆ �s��>�[���t6e{�b_'Q5F����!���"�^z�{�0����E_{����|��ʜ�]+�I�:hS���;~��DQ�<�*�T�d�Pe3Ӌ��y��^^��:A.�a.��{��5��k�6)ء3ӟ��ט��7���C����=�FD(
I�k��?U"ou����R<��S��0��"��ę��=��^E�cwƏU��d�����<��c0�K�ƾpT~�Cg4�ɂ�����}բ��Z��oא��ؿ��sF`~�4wm�����<�]�@�nhL�˗Z�GZ�3��b3gb��/|�wyZ��^�2�U���{�C�4��Z�y�,�tb2/�u��?4/*�PjW8W�t�噛Kwk�'��K������ň.Mt5��s]��j� ���B��E�Z1�əsf�tjA�:���۬�b����.���`���$}��aӕ��JWHA����@���A��OA��vy@q﵃յ���qX���c��D��Z:���a�<#x��t9i���Hv�Rq�a=��+k0%�:�n*��x#M�Z��_urvf9���Ʃy�l�3��1�J^��7�[�8��by�B3Z����t�\�����W�Z�[B�=�N�3c �U��f��=2p&v{�$�b�C&M���²q�c����>��>fL&ڱ9}򯷩���+�[� �t%e�.;�=
㎋#TT<�.��g�T%��C�%���!3�!@���,	Za�ͻ��m���n��r��Pd����7����cb�4�^���I��@��9�s<�Ryw���K�AJׄHR�C�mI� �|=��3�z�Ь�`����~Z���~�)�
:};0�݈�k�޻S��� ��CZ�b"�l&*�}`�B���$-�F���B��Dskrf��έ����tf�Z-DYh��T�j�}��F�$"��T-Os�e���$��R]�zJ�N43%��<T����dA}�E�D!y�>A����$;w�/�~80�=ٞ*��I��Ţ瓃��@���/����3�ޕ��&��;�����C��N�@�v���(<q�H�\4/K�<�1�xpF�ʭ�O� ��L`Y%�Q,=�k�*@����>�ʹI)Gv	gGw޻�l���(" ds�Y��{�]:{ߛ�&�
)t*�)���!����W�A��>}Ҵ�n͕N�.���8Y������-�ID��[�jY��f��	�b�Ơb)\@������EJ�n�v~m�]��iJՂ�LP��q���e�]5A7�TT��rQB�D�)Ĩ5C>��R�5�8��e�##�Tu=��߹+����<7��<y{��2)�
ʍ#��9U)e|��aG<�(*�I�:|�p��R^f�A�dޥ���΁gmK�2��ӹ�y��ߍL�������\��6y���R��Lfn��Ց[���g W��bs�}4�뫨�����`�~b�R����bgѭC6�Z3#�f�I$|��CB����F��{��y����N*Ƕ{Q�s��{Ε;�>�=�|�k�{6��Zx�]εA]��u�S���$\Na�*^���]�$��<ׅ_FwJZ���6���4:�u��C��s�_v(��'�w�[CՂ/&�<���J���_&Ǯ3":���1�����*��i�Ii
	����	͇(�t���V�}y�=G�� ��M�A��nz��wH��m���<#6�
������4A2����هB}�g�c����6��@��.�*�����A����n�E׽���O�6n ��LAˏ����~z�ׁ?��� ���*P%�&�3���w*O
�ø=�لp�ȁƺ@�}�+�:Y�}�su�6���7�!���R���*����ҮNJ&TI��-�73�u7��7S��?ʧp��cکg�CATH3��&F���:7�+}>��4^��~L-���wP�B��������âu���S�!оgI���~-�CtI�T��h�Vͭ������r��C̲��d��;�c~���L�$ä%��{��z��U觛We~���7�	��iE�0|�����	kûUц�2U6P��vq�e]�0���a?i�
Ċ��v	V],���="#�d�<\�Ⱥ�e�p�9֟v
<�*O��1C����|��~�䬡W��\4�پZS;�w��G�Ca�Uʰχ�n���>/��=w��G�N�%�|�.:���Q�Z�o����7�������4�D�$��˥������*��q�@���hFy�-�'r���C%����J����؋��-$Gu��))�����G���oe^G;:���>�=Yr5�b�T/_b�:�4'7�����Q�����v�S�/p�̹���t=2����P ��3�z}ԦˍNn��U!V�<���|�Pa�5��,�T��X��Lݍ��������Uy5�����+a�m��Z��T09�4�F�b|���jI�
���X�D�5�ƻhe]�dV�M����M�ڽ�>gޛz����fQ$�*�v�b���o��%`���Q�i$��/|�Ÿ5�΍;�U!�w�ɕ�5א���O�Uʐ��P�,-C1Gg�Ife��l�߲T�m��a��'Y5/k������͋=���8:�B���S�TB�Z2�����i����tQQ H*&9&"" �@I=
�˸d�o�4�ҡ>y�;&��VY�A�D��&2]
�]Ѭ�R��I�D)I�� ��R`�I D� �`�I�	�!Q���@�- " ��y �=9h�n��%�YB!�#��d�aH�EH� Q��9��i��煽F���ls�cP��W�o��>:��_��nߍGD�>�<3f������ �v��?Xvk�_,�._W}�>�`W �������aӠ<d=�b* ?$�!�*h^�3lov��C�0���S����}�4�Q���T ��8���ܹ"�HhÍ:ݠP 2��f�h�np��/ѿ��
K#7]k�W�_%3���T
��� � ���{�!�8�,�t% (B�CF�R�F-�o��KN����ٍ�l���j_^�P u�Bd7t��Q��iOv�<��R 3�
��,�@��q��oSX=�G����Y�����P! j�$p(<��U�[��s�Z���V�8h��8Cߵ��ِy�m�Yط/P���{2�g��j1�й� 0m�,������\9���.�Ѐ <U ߵ�F���/(����\�hN��&B�I �T��f䮸� �\��&5¨*��=�57�$���j�H>���d1��'3YJ%_-�J@�����P�X^���Q"v/Y�P d�� ��H�pP���j����)�ٳ�=��ң �S}&8�Ѱ0�ՈE:@�`C�I�w�=���(TD sh�y}*�0'o2�T �����c�/8fr�(�0mOU��M
^��r����[�P "�3�x��j�p����C;�-�cQ�[�̖o���+�re��ި 87�M)��s.���H�J�d�oE�\@ߎ���d1ŌI���.X\!��M@�h{J2Tw@�w]yl�����$~��!6��]�D� ��$�3�!vt����"�(HIw{�