BZh91AY&SY�%r� n_�Py����߰����`� x 1� @ @ " ��*�$��D�&F������A���(�   � ID�0�F ɂ�� �`�2��jy�Q$� H      `�1 �&	�!��L��IIO�M2�M�  ɚ'��pPR~�
"�� � ��}�,�+���wݨe�Ȁ��y켒��K�"���	�QD��g�ѳ �$dd�	E�$HEđ�	�	 	1I $		cFDd�@BD!EdXE �I�BEAR0	�! �	 $B@�	�%ӧ>?ꂽ��g�{��u��_��g�淗�����*j��ĀU�μҚ�ǌ�i�2ڳ]e��:;E4� �mTZh;fS&Êc:j6����ѡ����b�j�Қ#sd�c[+eqMGksv�����g��#�[P.�A�.����Wt�6`V`�LB�6\��
�[rF�0���k�)��h�L�,&,3�\��8ƷYenZ�;M�����l�*�Ö�j�[�,����Y�͚��XK��V��Z��R�h����5�9Ű�e��?n�-�{���K�t��x�G���պ�͟���v�8�3v^�w ���ш�B@&�*� �$dI�IX~I}�p�4! �Ʉ�;T1��v�+>����pܝ��<k��B,��:�r8㴮��ƺ��0a�]b@��G�̱���Μ�X���:�����<��0�_�6����$�1j�@B�DX�꠵�dӡ��$I���T�C�R����ӗ�_�U�٦w4`^��'i�0����^Qb&\x�>�*�<�<�73�""�LiXI��(!l�Đ�N
B�HL��� �J	/�*!�,䮙��8.�b���OA@`���ʏ���� �?���n�=�M/�@��8�08��*[b��A<����ٌfBm*~��Z��9�\��n��	K���DMD�\��>!�˻�>�$����	0ĖF�Tx�@25�T���U�9��?4{���k�� ��Y���2�BP��Cj({�|9�h�$��?t����T� � ZHÜo(Kn�+)Y�Ϫ��؄�@D"B��"� �9�ye�z(/Oe�����*�
��6�^ f�L\f	 6,k�u x;]q�ڄif�XFR�KZWn=/�<���݀�Z۫a5�I�O�B��AI�b���ˤ�I���m"����$s��H���'Ϙc��$�K~���lY�6|&V
�:�@T�Vg�w^%==�ZA�a�0چ!� �4x�w�SP�H�fQ.=e�4�P�阒7��`�a�/�
1���p�0����p���f�# vsA�25e�գ��C@���}y	VX�@X}��/j�9���K�m��ղ|&�}JEvȀ9�x�"�2�&�H��#�å'�;�"B������#9��0X�.���y4ʈ�L�� ���qE�a�6s.@v$6ts!��Ӊʠec�r�Di���#��%��)�����Vp���H1���pz:��P������j�V	�;�.�9{6���E@��}�\7yF��Z�$���u�R�y��mi�P�Q�����mв�����4��Ҧ͋��� �.0��^��lbt"�vxb�bff^���w�rBf
���U��`�+#6�Q#�	��>4�.�l�.�����Aż-�,���@,"�p@O��N�qc��־!`Zƃ�vzN�Ҷ�b��ب�\^d�ʀ���f��|eB�L&��a�r�#���pH�62�^���e���i�yX����IuS]@�ѳFjh�0~7��0�-&� $\@P+� ���M�
��.Ø,���I����pY	�t1���t�WR3Պn���zKV��K�!؍b� �,��yTů�s�0��W�O�C�zyn��v^�I�;]t���l�2��u�m�m�CM��[2�2b1[���&e�H�7+-n^�ERB."|De��n�����+�H��������Ͱ�R����]\j�I��v22��MDJŉQ� �E���,�����B;�/Q�:䊻$�q1� �/n62&���݈���F�9��=
 C>P� ��Q"�T���wm�Ӻ+���$Q�,���Ω����ݽ�\`�݃L�K�jȌ�h��"(��!��N���`N+��Bh�|;�E���x����]��� �֐RVq٦�*;`I���(�n#|F.~���PC(c^�\'J�v �����B�@�uK�gtH� �f�+sn�i�K�i[�5�c����Z:���tj$�� �abK��l�a@��L���/�����I�m�*���B$�Q�3�>JEA��6��8[�\u����n(�ۜ���}�Wj\��,+r�E���H�y�+�3fS�}sS�()/"Ve����/9����<Y�Nʋ��<uY�s4��f@mD$"!��
i�8p�c�#n�&�G@�u�\�=���k��G��)�;7MH����np%A�J &�F[��ד)wU�e�F[٦�%f0J5��Kr�o��%{�\��h��d��Y
�E���z��A�u,�k�1{b(R�$ir!pg�d�e�]C�ĉ�R7�����$!'�I$�
QG�@����	��(��k���v�����X�a�-�
 �E4Zb�QKK�J�HAL��j)kB�(���0����]���~VueZ�J$5�����c�@BID�ʧ�k9;9Gy)짿q�0���Q�|���m�\�&��� ���$}�4�q3ͧש��!��RǦ�\\Prq�����	���V�!֊�m�7Q=��4;S��,�w��]{�B�������!��D��t���/<w��2vg�dzN ,L���L!���0��q��^ QAYe����f�q������ZD��4�X�mF��R� vDA@D��%U4ذ]�X�YƭE��,`n�Ԝ?�Xd�� Me.pl�֑�A�9�&Ҍ�j04lC2�RFp�V|{�A���.zƻ'E��qy�h�E@S"�I��ry��x|S��=<��
^m�5X1ٰĸ�9�S#�@:���ܩ�A�aE�C� �Zف�!����v]�Npc� ���M�: )�o}B@7�1�f��M�&��+~Tmt&�Ũ��j6�`2���\	�l�Q� ���p�Gqǀ,�h�v�(�~%<v#�4�NyQ�ސ�&;Ӄ��&R�pH8&���� J�耧ؠ>�$~�3�܆�k,<���o�3)7�v�ͪ#�
����6Й�R�*[�<��7G��~�g0������X�# �<�Έ
d6>�;��}f��Pr�7���mC2G4h�����Y\i�!RĘv9'���/Ub��L�P� �Q�b*&�sV�l"��@1�n6`�EQ�nl�d�?�K��B�{kh�5���#���!vs��6E>IGYf��,���ä7�m����I�T��1"Y��/�W!	�J������rE8P��%r�